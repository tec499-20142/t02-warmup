module warmup(
	input wire clk,
	input wire rsPin);

	uart rs232();
	
	always @(posedge clk)
		begin
		
		end
endmodule